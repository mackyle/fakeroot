PO4A-HEADER:mode=after;position=FÖRFATTARE;beginboundary=.SH
.SH ÖVERSÄTTNING
David Weinehall
.RI < tao@kernel.org >
